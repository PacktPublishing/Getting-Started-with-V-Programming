module mod1

const greet_count = 5

pub fn do_work() {
	println(mod1.greet_count)
}
