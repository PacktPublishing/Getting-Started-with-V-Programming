module main

fn main() {
	a := 10
	b := 2

	// add using +
	sum := a + b

	// subtract using -
	diff := b - a

	// product using *
	prod := a * b

	// / results in quotient
	quotient := a / b

	// % modulo results in remainder
	remainder := a % b

	println('Sum of $a and $b is $sum')
	println('Subtracting $a from $b is $diff')
	println('Product of $a and $b is $prod')
	println('Quotient when $a divided by $b is $quotient')
	println('Remainder when $a divided by $b is $remainder')
}
