module main

fn main() {
	i := 'hello' // i is not used anywhere, so warns when run in dev mode and throws error when run in prod mode
	x := 3
	y := 2
	println(x + y)
}
