module main

import m1
import m2

fn main() {
	m1.hello()
	m2.hello()
}
