module main

fn method1() {
	msg := 'Hello from Method1'
	println(msg)
}

fn method2() {
	msg := 'Hello from Method2'
	println(msg)
}

fn main() {
	method1()
	method2()
}
