module mod1

pub fn hello2() {
	println('Hello 2 from mod1!')
}
