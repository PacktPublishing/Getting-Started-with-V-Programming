module mod1

pub fn hello() string {
	return 'Hello from mod1!'
}
