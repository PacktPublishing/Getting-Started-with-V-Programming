module mod1

pub fn hello() {
	println('Hello from mod1!')
}
