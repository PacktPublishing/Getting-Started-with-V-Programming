module main

fn main() {
	println('Welcome to the World of V!')
}
