module mod1

pub const greet_msg = 'Greeting from mod1!'
