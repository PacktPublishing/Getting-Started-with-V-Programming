module main

import mod1

fn main() {
	println(mod1.greet_msg)
}
