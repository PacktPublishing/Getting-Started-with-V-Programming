module main

import mod1

fn main() {
	println('Hello World!')
}
