module main

// greet function prints greetings to the console
pub fn greet() {
	println('Hello, Welcome to the Jungle!')
}

fn main() {
	greet()
}
