module main

fn main() {
        hs := 'Monday'

        if hs.contains('mon') {
                println('$hs contains mon')
        } else {
                println('$hs does not contains mon')
        }
}
