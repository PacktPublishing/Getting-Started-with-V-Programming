module main

const app_name = 'V on Wheels'

fn main() {
	println(app_name)
}
