module mod1

pub fn hello() {
	println('Hello from mod1!')
}

fn init() {
	println('Initializing mod1')
}
