module main

fn main() {
	hs := 'monday'

	if hs.contains('mon') {
		println('$hs contains mon')
	} else {
		println('$hs does not contains mon')
	}
}
