module main

import mod1

fn main() {
	mod1.hello()
	println('Hello World!')
}
