module mod1

fn hello2() {
	println('Hello 2 from mod1!')
}
