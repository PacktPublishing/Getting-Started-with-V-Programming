module main

import mod1

fn main() {
	res := mod1.hello()
	println(res)
}
