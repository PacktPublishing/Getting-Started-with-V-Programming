module main

import mod1

fn main() {
	mod1.do_work()
}
