// file: mymod/mymod.v
module mymod

__global (
	msg string
)
